module InstMem (input [5:0] addr, output [31:0] data_out);
reg [31:0] mem [0:63];
initial begin

mem[0]  = 32'b00000000111100000000000110010011; 
mem[1]  = 32'b00000001010000000000000010010011;
mem[2]  = 32'b00000010010000001000000100010011; 
mem[3]  = 32'b00000000001100010000000010110011;
mem[4]  = 32'b01000000001100010000000010110011;
mem[5]  = 32'b00000000001100010100000010110011;
mem[6]  = 32'b00000000001100010110000010110011;
mem[7]  = 32'b00000000001100010111000010110011;
mem[8]  = 32'b00000000001100010001000010110011;
mem[9]  = 32'b00000000001100010101000010110011;
mem[10] = 32'b01000000001100010101000010110011;
mem[11] = 32'b00000000001100010010000010110011;
mem[12] = 32'b00000000001100010011000010110011;
mem[13] = 32'b00000000001000010000000010010011;
mem[14] = 32'b00000000001000010100000010010011;
mem[15] = 32'b00000000001000010110000010010011;
mem[16] = 32'b00000000001000010111000010010011;
mem[17] = 32'b00000000001000010001000010010011;
mem[18] = 32'b00000000001100010101000010010011;
mem[19] = 32'b01000000001100010101000010010011;
mem[20] = 32'b00000000001100010010000010010011;
mem[21] = 32'b00000000001100010011000010010011;
mem[22] = 32'b00000000000100010000000100100011; //sb
mem[23] = 32'b00000000000100010001000100100011;
mem[24] = 32'b00000000000100010010000100100011;
mem[25] = 32'b00000000001000010000000010000011;
mem[26] = 32'b00000000001000010001000010000011;
mem[27] = 32'b00000000001000010010000010000011;
mem[28] = 32'b00000000001000010100000010000011;
mem[29] = 32'b00000000001000010101000010000011; 
mem[30] = 32'b00000000001000001000001001100011;
mem[31] = 32'b00000000001000001001001001100011;
mem[32] = 32'b00000000001000001100001001100011;
mem[33] = 32'b00000000001000001101001001100011;
mem[34] = 32'b00000000001000001110001001100011;
mem[35] = 32'b00000000001000001111001001100011;
mem[36] = 32'b00000000000000001100000010110111;
mem[37] = 32'b00000000000000001100000010010111;
mem[38] = 32'b00000000000000000000000001110011;

end
assign data_out = mem[addr];

endmodule